module hex_to_binary (
    input  [15:0] H,     // 16 one-hot inputs
    output reg [3:0] B   // 4-bit binary output
);
always @(*) begin
    case (H)
        16'b0000000000000001: B = 4'b0000; // 0
        16'b0000000000000010: B = 4'b0001; // 1
        16'b0000000000000100: B = 4'b0010; // 2
        16'b0000000000001000: B = 4'b0011; // 3
        16'b0000000000010000: B = 4'b0100; // 4
        16'b0000000000100000: B = 4'b0101; // 5
        16'b0000000001000000: B = 4'b0110; // 6
        16'b0000000010000000: B = 4'b0111; // 7
        16'b0000000100000000: B = 4'b1000; // 8
        16'b0000001000000000: B = 4'b1001; // 9
        16'b0000010000000000: B = 4'b1010; // A
        16'b0000100000000000: B = 4'b1011; // B
        16'b0001000000000000: B = 4'b1100; // C
        16'b0010000000000000: B = 4'b1101; // D
        16'b0100000000000000: B = 4'b1110; // E
        16'b1000000000000000: B = 4'b1111; // F
        default: B = 4'b0000; // Invalid input
    endcase
end
